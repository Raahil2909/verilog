`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:59:03 01/19/2021 
// Design Name: 
// Module Name:    carrry_look_ahead 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module carrry_look_ahead(
    input [3:0] a,
    input [3:0] b,
    input c,
    output [3:0] s,
    output cout
    );
wire p0,p1,p2,p3,g0,g1,g2,g3,c1,c2,c3,c4;

assign #2 p0=(a[0]^b[0]),
       p1=(a[1]^b[1]),
       p2=(a[2]^b[2]),
       p3=(a[3]^b[3]);
		 
assign #2 g0=(a[0]&b[0]),
       g1=(a[1]&b[1]),
       g2=(a[2]&b[2]),
       g3=(a[3]&b[3]);
		 
assign #2 c0=c,
       c1=g0|(p0&c),
       c2=g1|(p1&g0)|(p1&p0&c),
       c3=g2|(p2&g1)|(p2&p1&g0)|(p1&p1&p0&c),
       c4=g3|(p3&g2)|(p3&p2&g1)|(p3&p2&p1&g0)|(p3&p2&p1&p0&c);
		 
assign #2 s[0]=p0^c0,
       s[1]=p1^c1,
       s[2]=p2^c2,
       s[3]=p3^c3;
		 
assign cout=c4;

endmodule
